`ifndef DUV_TYPE_GUARD
`define DUV_TYPE_GUARD
	typedef enum logic { SIN_SEGMENTAR, SEGMENTADO } e_duv_type;
`endif